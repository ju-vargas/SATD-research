`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:01:19 10/27/2023 
// Design Name: 
// Module Name:    SATD_tb 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 

//////////////////////////////////////////////////////////////////////////////////
module SATD_tb(
    );

	//parametros
   parameter CLK_PERIOD = 2;  
	integer count = 0;
	//sinais de testbench
	reg clk;
	reg reset;
	
	//entradas e saidas pra teste
	wire [1023:0] input_ORG; 
	wire [1023:0] input_CUR;
	
	
	//module instantiation 		
	SATD #( .WIDTH (8), .NUM_INPUTS (8), .ITERATIONS (15)) satd
	       (	.clk 	 		  	(clk),
				.rst	 		  	(reset),
				.ORG 			  	(input_ORG),
				.CUR 			  	(input_CUR));
					
    //NUM_INPUTS !!SEMPRE 8!!, por enquanto
    //  --pq eu nao consigo mudar o numero de registradores q to usando. 
	//assign input_ORG = {60'b0, 4'b1111};
	//assign input_CUR = {60'b0, 4'b0011};
	
	assign input_ORG = {64'b0011011010101101111010110011001100110011001110111101101101001001,
							  64'b0101010101010101010101010101010101010101010101010101010101010101,
							  64'b0011001100110011001100110011001100110011001100110011001100110011,
							  64'b1100110011001100110011001100110011001100110011001100110011001100,
							  64'b0000111100001111000011110000111100001111000011110000111100001111,
							  64'b1111000011110000111100001111000011110000111100001111000011110000,
							  64'b0100010001000100010001000100010001000100010001000100010001000100,
							  64'b1001111111111111111110001000100010001000100010001000100010001000,
							  64'b0000000000000000000000000111111110000000011111111000000001111111,
							  64'b1111111100000000111111110000000011111111000000001111111000000000,
							  64'b0101010010101010101010101010010101010101010101010101010101010101,
							  64'b1010101001010101010101010101101010101010101010101010101010101101,
							  64'b1100110011110011001100110011110011001100110011110011001100110011,
							  64'b0011001100001100110011001100001100110011001100001100110011001100,
							  64'b0000111100001111000011110000111100001111000011110000111100011111,
							  64'b1111000011110000111100001111000111100001111000111100001111110000};
					
					
	assign input_CUR = {64'b1011001001011110100101100110000010011001000111111001101000111111,
							  64'b1111110101010101010101010101010101010101010101010101010101010101,
							  64'b1011001100011010101100111100110001101001111001001111001001000110,
							  64'b0011111000110111001000110011001011111100011101001111110101100100,
							  64'b0101010101010100011100010100011101010011001010001010000101000100,
							  64'b1111000011000000111101010000100011111001101001010101000000000010,
							  64'b0100000100101000100001000101000010001010001001000100010000000000,
							  64'b1000010010010001001000100001000100010001000010010001000100000000,
							  64'b0000000011111111100000000111111110000000011111111000000001111111,
							  64'b1111111000000000000011111111000000000000011111110000000000000000,
							  64'b0010001000101010101010010101001001010000101010101001001010010101,
							  64'b1001010100010101001001010101001101000101010101010101010001000101,
							  64'b1111010011110111001100110011110011010101111010011001110001001100,
							  64'b1111111111111111111111111111111111111111111111111110011001100110,
							  64'b0100011000100010001010010101000010001001000101000001001000010001,
							  64'b1111111111111111111111111111111111111111010001010101000101010101};
									  
	initial begin
		clk   <= 0;
		reset <= 1;
	end
	
	//geracao do sinais		
	always begin
		#CLK_PERIOD clk = ~clk; 
		  
		reset <= 0;

      count = count + 1;
      if (count == CLK_PERIOD*30) begin
          $stop; 
		end	
	end

endmodule
